// hello.v
module hello;
  initial begin
    $display("Hello from Verilator!");
    $finish;
  end
endmodule
