module TopModule();

  
endmodule
