module TopModule();
endmodule
