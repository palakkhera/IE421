/*
BRAM --> Block Random Access Memory
  Used to store large amounts of memory in your FPGA
  Close proximity to the FPGA logic circuits --> high speed access 
  Good for rapid retrieval 
  Often used to store Lookup tables

Inputs:
Outputs:
Goal:
  Implement a True Dual Port BRAM
  Provide fast and effienct memory storage for data and intructions
*/

module bram (input logic variable_in
             output logic variable_out);
endmodule

